module JKflipflop (
    input j,k,clk, output reg q, output qbar      // this is when assign statement is used, maybe ok 
    // inout j,k,clk, output reg q,qbar
);

    always @(posedge clk) begin
        q <= (j& ~q) | (~k & q);
        
    end
    assign qbar = ~q;

    // always @(posedge clk) begin             // this is purely sequential circuit
    //     case({j,k})
    //         2'b00: begin q<=q; qbar<=qbar; end
    //         2'b01: begin q<=1'b0; qbar<=1'b1; end
    //         2'b10: begin q<=1'b1; qbar<=1'b0; end
    //         2'b11: begin q<= ~q; qbar<= ~qbar; end
    //         default : q<=x; qbar<=x;
    //     endcase    
    // end
            
endmodule
